module main

fn main() {
	println('Hello, World!')
}

fn greet(name string) string {
	return 'Hello, ${name}!'
}